module od_buf(y, a);
	input wire a;
	output wire y;
	
	assign y = a;

endmodule